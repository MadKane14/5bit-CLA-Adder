* SPICE3 file created from inverter.ext - technology: scmos
.include TSMC_180nm.txt

Vdd Vdd 0 1.8
Vin IN 0 PULSE(0 1.8 0 0n 0n 1n 2n)

M1000 OUT IN Vdd Vdd CMOSP w=1.8u l=0.18u
M1001 OUT IN 0   0   CMOSN w=0.9u l=0.18u

C0 IN Vdd 0.06fF
C1 OUT Vdd 0.28fF
C2 0 OUT 0.13fF
C3 IN OUT 0.05fF
C4 0 0 0.17fF
C5 OUT 0 0.10fF
C6 IN 0 0.22fF
C7 Vdd 0 1.21fF

.tran 0.1n 10n

.control
set color0 = white
set color1 = black

run
set curplottitle="Madhur-Kankane-2024102061-3-OR"
plot V(IN) 2+V(OUT)

.endc
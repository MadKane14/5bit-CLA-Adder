* SPICE3 file created from and.ext - technology: scmos
.include TSMC_180nm.txt

Vdd Vdd 0 1.8
Va a 0 PULSE(0 1.8 0 0n 0n 5n 10n)
Vb b 0 PULSE(0 1.8 0 0n 0n 10n 20n)

M1000 y nand_0/y Vdd Vdd CMOSP w=1.8u l=0.18u
M1001 y nand_0/y 0   0   CMOSN w=0.9u l=0.18u

M1002 Vdd a nand_0/y Vdd CMOSP w=1.8u l=0.18u
M1005 nand_0/y b Vdd Vdd CMOSP w=1.8u l=0.18u


M1004 nand_0/y a nand_0/a_57_n34# 0 CMOSN w=0.9u l=0.18u
M1003 nand_0/a_57_n34# b 0 0 CMOSN w=0.9u l=0.18u

C0 a Vdd 0.06fF
C1 b Vdd 0.06fF
C2 b a 0.42fF
C3 b 0 0.04fF
C4 y Vdd 0.28fF
C5 y 0 0.13fF
C6 nand_0/y Vdd 0.48fF
C7 nand_0/y a 0.23fF
C8 nand_0/y 0 0.03fF
C9 nand_0/y y 0.05fF
C10 Vdd 0 3.00fF
C11 a 0 0.26fF
C12 b 0 0.24fF
C13 0 0 0.31fF
C14 y 0 0.12fF
C15 nand_0/y 0 0.35fF

.tran 0.1n 40n

.control
set color0 = white
set color1 = black

run
set curplottitle="Madhur-Kankane-2024102061-3-AND"
plot V(a) 2+V(b) 4+V(y)

.endc

* SPICE3 file created from or.ext - technology: scmos
.include TSMC_180nm.txt

Vdd Vdd 0 1.8
Va a 0 PULSE(0 1.8 0 0n 0n 5n 10n)
Vb b 0 PULSE(0 1.8 0 0n 0n 10n 20n)


M1000 y nor_0/y Vdd Vdd CMOSP w=1.8u l=0.18u
M1001 y nor_0/y 0   0   CMOSN w=0.9u l=0.18u

M1002 nor_0/a_65_6# b Vdd Vdd CMOSP w=1.8u l=0.18u
M1005 nor_0/y a nor_0/a_65_6# Vdd CMOSP w=1.8u l=0.18u

M1003 nor_0/y b 0 0 CMOSN w=0.9u l=0.18u
M1004 0 a nor_0/y 0 CMOSN w=0.9u l=0.18u

C0 a b 0.43fF
C1 nor_0/y a 0.13fF
C2 Vdd b 0.06fF
C3 Vdd a 0.06fF
C4 Vdd nor_0/y 0.09fF
C5 nor_0/y 0 0.21fF
C6 y nor_0/y 0.05fF
C7 Vdd y 0.28fF
C8 y 0 0.13fF
C9 Vdd 0 3.05fF
C10 0 0 0.34fF
C11 nor_0/y 0 0.36fF
C12 a 0 0.26fF
C13 b 0 0.24fF
C14 y 0 0.13fF

.tran 0.1n 40n

.control
set color0 = white
set color1 = black

run
set curplottitle="Madhur-Kankane-2024102061-6-OR"
plot V(a) 2+V(b) 4+V(y)

.endc